--------------------------------------------------------------------------------
-- PIA
-- THIEBOLT Francois Janvier 2014
--------------------------------------------------------------------------------

-- Definition des librairies
library IEEE;
library STD;

-- Definition des portee d'utilisation
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use IEEE.std_logic_unsigned.all;

-- -----------------------------------------------------------------------------
-- Definition de l'entite
-- -----------------------------------------------------------------------------
entity pia is

	-- definition des parametres generiques
  generic	(
		-- largeur par defaut des bus
    IOSIZE : ________ );

	-- definition des entrees/sorties
  port 	(
		-- signaux de controle du cache
		___________
		___________
		___________
		___________
		___________ );

end pia;


-- -----------------------------------------------------------------------------
-- Definition de l'architecture du pia
-- -----------------------------------------------------------------------------
architecture behavior of pia is

	-- definition de constantes

	-- declaration des ressources locales
	___________
	___________
	___________


begin
--------------------------------------------
-- Affectations dans le domaine combinatoire
_________
_________
_________
_________

---------------------
-- Process PIA ACCESS
PIA_ACCESS: process(__________)
begin
	___________
	___________
	___________
	___________
	___________
	___________
	___________
	___________
	___________
	___________
	___________
	___________
	___________
	___________
	___________

end process PIA_ACCESS;

end behavior;

